//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module add
(
  input  [3:0] a, b,
  output [3:0] sum
);

  assign sum = a + b;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module signed_add_with_overflow
(
  input  [3:0] a, b,
  output [3:0] sum,
  output     logic  overflow
);
  
    add a1 (.a(a)    ,
            .b(b)    ,
            .sum(sum));
  
    assign overflow = ((a[3] & b[3] & ~sum[3]) || (~a[3] & ~b[3] & sum[3]));

endmodule
