//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux
(
  input  d0, d1,
  input  sel,
  output y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module not_gate_using_mux
(
    input  i,
    output o
);

wire z = 0;
wire x = 1;

mux m (
  .d0 (x),
  .d1 (z), 
  .sel (i),
  .y (o)
  );

endmodule
