//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux
(
  input  d0, d1,
  input  sel,
  output y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module xor_gate_using_mux
(
    input  a,
    input  b,
    output o
);

wire z = 0;
wire x = 1;
wire b_n;

mux n (
  .d0 (x),
  .d1 (z), 
  .sel (b),
  .y (b_n)
  );

mux m (
  .d0 (b),
  .d1 (b_n), 
  .sel (a), 
  .y (o)
  ); 



endmodule
